`timescale 1ns / 1ps

module testbench();
    reg [3:0] d1, d0, sh_amt;
    reg sel, clk, rst;
    wire gt, lt, eq;
    wire [3:0] regOut, sum, diff, prod, muxOut, shrOut, shlOut, quot, rem, incOut, decOut;
    
    REG #(.DATAWIDTH(4)) reg1(d0, regOut, clk, rst);
    ADD #(.DATAWIDTH(4)) add1(d1,d0,sum);
    SUB #(.DATAWIDTH(4)) sub1(d1,d0,diff);
    MUL #(.DATAWIDTH(4)) mul1(d1,d0,prod);
    COMP #(.DATAWIDTH(4)) comp(d1,d0,gt,lt,eq);
    MUX2x1 #(.DATAWIDTH(4)) mux1(d1,d0,sel,muxOut);
    SHR #(.DATAWIDTH(4)) shr1(d0,sh_amt,shrOut);
    SHL #(.DATAWIDTH(4)) shl1(d0,sh_amt,shlOut);
    DIV #(.DATAWIDTH(4)) div1(d1,d0,quot);
    MOD #(.DATAWIDTH(4)) mod1(d1,d0,rem);
    INC #(.DATAWIDTH(4)) inc1(d0,incOut);
    DEC #(.DATAWIDTH(4)) dec1(d0,decOut);
    
    initial begin
        clk <= 0;
        #10 rst <= 0; sh_amt = 0; d1 <= 0; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 0; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 0; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 0; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 0; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 0; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 0; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 0; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 0; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 0; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 0; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 0; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 0; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 0; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 0; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 0; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 0; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 0; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 0; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 0; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 0; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 0; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 0; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 0; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 0; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 0; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 0; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 0; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 0; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 0; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 0; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 0; d0 <= 15; sel <= 1; // 
        #10 rst <= 0; sh_amt = 0; d1 <= 1; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 1; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 1; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 1; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 1; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 1; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 1; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 1; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 1; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 1; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 1; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 1; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 1; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 1; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 1; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 1; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 1; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 1; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 1; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 1; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 1; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 1; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 1; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 1; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 1; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 1; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 1; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 1; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 1; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 1; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 1; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 1; d0 <= 15; sel <= 1; // 
        #10 rst <= 0; sh_amt = 0; d1 <= 2; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 2; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 2; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 2; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 2; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 2; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 2; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 2; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 2; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 2; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 2; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 2; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 2; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 2; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 2; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 2; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 2; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 2; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 2; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 2; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 2; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 2; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 2; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 2; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 2; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 2; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 2; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 2; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 2; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 2; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 2; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 2; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 3; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 3; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 3; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 3; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 3; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 3; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 3; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 3; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 3; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 3; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 3; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 3; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 3; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 3; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 3; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 3; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 3; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 3; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 3; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 3; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 3; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 3; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 3; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 3; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 3; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 3; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 3; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 3; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 3; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 3; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 3; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 3; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 4; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 4; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 4; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 4; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 4; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 4; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 4; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 4; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 4; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 4; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 4; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 4; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 4; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 4; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 4; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 4; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 4; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 4; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 4; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 4; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 4; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 4; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 4; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 4; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 4; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 4; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 4; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 4; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 4; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 4; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 4; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 4; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 5; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 5; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 5; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 5; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 5; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 5; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 5; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 5; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 5; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 5; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 5; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 5; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 5; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 5; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 5; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 5; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 5; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 5; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 5; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 5; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 5; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 5; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 5; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 5; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 5; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 5; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 5; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 5; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 5; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 5; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 5; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 5; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 6; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 6; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 6; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 6; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 6; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 6; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 6; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 6; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 6; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 6; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 6; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 6; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 6; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 6; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 6; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 6; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 6; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 6; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 6; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 6; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 6; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 6; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 6; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 6; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 6; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 6; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 6; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 6; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 6; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 6; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 6; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 6; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 7; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 7; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 7; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 7; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 7; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 7; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 7; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 7; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 7; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 7; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 7; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 7; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 7; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 7; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 7; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 7; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 7; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 7; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 7; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 7; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 7; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 7; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 7; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 7; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 7; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 7; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 7; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 7; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 7; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 7; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 7; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 7; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 8; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 8; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 8; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 8; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 8; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 8; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 8; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 8; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 8; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 8; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 8; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 8; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 8; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 8; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 8; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 8; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 8; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 8; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 8; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 8; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 8; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 8; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 8; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 8; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 8; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 8; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 8; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 8; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 8; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 8; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 8; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 8; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 9; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 9; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 9; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 9; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 9; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 9; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 9; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 9; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 9; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 9; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 9; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 9; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 9; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 9; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 9; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 9; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 9; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 9; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 9; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 9; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 9; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 9; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 9; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 9; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 9; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 9; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 9; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 9; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 9; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 9; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 9; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 9; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 10; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 10; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 10; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 10; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 10; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 10; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 10; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 10; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 10; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 10; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 10; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 10; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 10; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 10; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 10; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 10; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 10; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 10; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 10; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 10; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 10; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 10; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 10; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 10; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 10; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 10; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 10; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 10; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 10; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 10; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 10; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 10; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 11; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 11; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 11; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 11; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 11; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 11; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 11; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 11; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 11; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 11; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 11; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 11; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 11; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 11; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 11; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 11; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 11; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 11; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 11; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 11; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 11; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 11; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 11; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 11; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 11; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 11; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 11; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 11; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 11; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 11; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 11; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 11; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 12; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 12; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 12; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 12; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 12; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 12; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 12; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 12; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 12; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 12; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 12; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 12; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 12; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 12; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 12; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 12; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 12; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 12; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 12; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 12; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 12; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 12; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 12; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 12; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 12; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 12; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 12; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 12; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 12; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 12; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 12; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 12; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 13; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 13; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 13; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 13; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 13; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 13; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 13; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 13; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 13; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 13; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 13; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 13; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 13; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 13; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 13; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 13; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 13; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 13; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 13; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 13; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 13; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 13; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 13; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 13; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 13; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 13; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 13; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 13; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 13; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 13; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 13; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 13; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 14; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 14; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 14; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 14; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 14; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 14; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 14; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 14; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 14; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 14; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 14; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 14; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 14; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 14; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 14; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 14; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 14; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 14; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 14; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 14; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 14; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 14; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 14; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 14; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 14; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 14; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 14; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 14; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 14; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 14; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 14; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 14; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 15; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 15; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 15; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 15; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 15; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 15; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 15; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 15; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 15; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 15; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 15; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 15; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 15; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 15; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 15; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 15; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 15; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 15; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 15; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 15; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 15; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 15; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 15; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 15; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 15; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 15; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 15; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 15; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 15; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 0; d1 <= 15; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 0; d1 <= 15; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 15; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 0; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 0; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 0; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 0; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 0; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 0; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 0; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 0; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 0; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 0; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 0; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 0; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 0; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 0; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 0; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 0; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 0; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 0; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 0; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 0; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 0; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 0; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 0; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 0; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 0; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 0; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 0; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 0; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 0; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 0; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 0; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 0; d0 <= 15; sel <= 1; // 
        #10 rst <= 0; sh_amt = 1; d1 <= 1; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 1; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 1; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 1; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 1; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 1; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 1; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 1; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 1; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 1; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 1; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 1; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 1; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 1; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 1; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 1; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 1; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 1; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 1; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 1; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 1; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 1; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 1; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 1; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 1; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 1; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 1; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 1; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 1; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 1; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 1; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 1; d0 <= 15; sel <= 1; // 
        #10 rst <= 0; sh_amt = 1; d1 <= 2; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 2; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 2; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 2; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 2; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 2; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 2; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 2; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 2; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 2; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 2; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 2; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 2; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 2; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 2; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 2; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 2; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 2; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 2; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 2; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 2; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 2; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 2; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 2; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 2; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 2; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 2; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 2; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 2; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 2; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 2; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 2; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 3; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 3; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 3; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 3; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 3; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 3; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 3; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 3; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 3; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 3; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 3; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 3; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 3; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 3; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 3; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 3; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 3; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 3; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 3; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 3; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 3; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 3; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 3; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 3; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 3; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 3; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 3; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 3; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 3; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 3; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 3; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 3; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 4; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 4; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 4; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 4; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 4; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 4; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 4; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 4; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 4; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 4; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 4; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 4; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 4; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 4; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 4; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 4; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 4; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 4; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 4; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 4; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 4; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 4; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 4; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 4; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 4; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 4; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 4; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 4; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 4; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 4; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 4; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 4; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 5; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 5; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 5; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 5; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 5; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 5; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 5; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 5; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 5; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 5; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 5; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 5; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 5; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 5; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 5; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 5; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 5; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 5; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 5; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 5; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 5; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 5; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 5; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 5; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 5; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 5; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 5; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 5; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 5; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 5; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 5; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 5; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 6; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 6; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 6; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 6; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 6; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 6; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 6; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 6; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 6; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 6; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 6; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 6; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 6; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 6; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 6; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 6; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 6; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 6; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 6; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 6; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 6; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 6; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 6; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 6; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 6; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 6; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 6; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 6; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 6; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 6; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 6; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 6; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 7; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 7; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 7; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 7; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 7; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 7; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 7; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 7; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 7; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 7; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 7; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 7; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 7; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 7; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 7; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 7; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 7; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 7; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 7; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 7; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 7; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 7; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 7; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 7; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 7; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 7; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 7; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 7; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 7; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 7; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 7; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 7; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 8; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 8; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 8; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 8; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 8; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 8; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 8; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 8; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 8; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 8; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 8; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 8; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 8; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 8; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 8; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 8; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 8; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 8; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 8; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 8; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 8; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 8; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 8; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 8; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 8; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 8; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 8; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 8; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 8; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 8; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 8; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 8; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 9; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 9; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 9; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 9; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 9; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 9; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 9; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 9; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 9; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 9; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 9; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 9; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 9; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 9; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 9; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 9; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 9; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 9; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 9; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 9; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 9; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 9; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 9; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 9; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 9; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 9; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 9; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 9; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 9; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 9; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 9; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 9; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 10; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 10; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 10; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 10; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 10; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 10; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 10; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 10; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 10; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 10; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 10; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 10; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 10; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 10; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 10; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 10; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 10; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 10; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 10; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 10; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 10; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 10; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 10; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 10; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 10; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 10; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 10; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 10; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 10; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 10; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 10; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 10; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 11; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 11; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 11; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 11; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 11; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 11; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 11; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 11; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 11; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 11; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 11; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 11; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 11; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 11; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 11; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 11; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 11; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 11; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 11; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 11; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 11; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 11; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 11; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 11; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 11; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 11; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 11; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 11; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 11; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 11; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 11; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 11; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 12; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 12; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 12; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 12; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 12; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 12; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 12; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 12; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 12; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 12; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 12; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 12; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 12; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 12; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 12; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 12; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 12; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 12; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 12; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 12; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 12; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 12; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 12; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 12; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 12; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 12; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 12; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 12; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 12; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 12; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 12; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 12; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 13; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 13; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 13; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 13; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 13; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 13; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 13; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 13; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 13; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 13; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 13; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 13; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 13; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 13; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 13; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 13; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 13; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 13; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 13; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 13; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 13; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 13; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 13; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 13; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 13; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 13; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 13; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 13; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 13; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 13; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 13; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 13; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 14; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 14; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 14; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 14; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 14; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 14; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 14; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 14; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 14; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 14; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 14; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 14; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 14; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 14; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 14; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 14; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 14; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 14; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 14; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 14; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 14; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 14; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 14; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 14; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 14; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 14; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 14; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 14; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 14; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 14; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 14; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 14; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 15; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 15; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 15; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 15; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 15; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 15; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 15; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 15; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 15; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 15; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 15; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 15; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 15; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 15; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 15; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 15; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 15; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 15; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 15; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 15; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 15; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 15; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 15; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 15; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 15; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 15; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 15; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 15; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 15; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 15; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 1; d1 <= 15; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 1; d1 <= 15; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 0; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 0; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 0; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 0; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 0; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 0; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 0; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 0; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 0; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 0; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 0; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 0; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 0; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 0; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 0; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 0; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 0; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 0; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 0; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 0; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 0; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 0; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 0; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 0; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 0; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 0; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 0; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 0; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 0; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 0; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 0; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 0; d0 <= 15; sel <= 1; // 
        #10 rst <= 0; sh_amt = 2; d1 <= 1; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 1; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 1; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 1; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 1; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 1; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 1; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 1; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 1; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 1; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 1; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 1; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 1; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 1; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 1; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 1; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 1; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 1; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 1; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 1; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 1; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 1; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 1; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 1; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 1; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 1; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 1; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 1; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 1; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 1; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 1; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 1; d0 <= 15; sel <= 1; // 
        #10 rst <= 0; sh_amt = 2; d1 <= 2; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 2; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 2; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 2; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 2; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 2; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 2; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 2; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 2; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 2; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 2; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 2; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 2; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 2; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 2; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 2; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 2; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 2; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 2; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 2; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 2; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 2; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 2; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 2; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 2; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 2; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 2; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 2; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 2; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 2; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 2; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 2; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 3; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 3; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 3; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 3; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 3; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 3; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 3; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 3; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 3; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 3; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 3; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 3; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 3; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 3; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 3; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 3; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 3; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 3; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 3; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 3; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 3; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 3; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 3; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 3; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 3; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 3; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 3; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 3; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 3; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 3; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 3; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 3; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 4; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 4; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 4; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 4; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 4; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 4; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 4; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 4; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 4; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 4; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 4; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 4; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 4; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 4; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 4; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 4; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 4; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 4; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 4; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 4; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 4; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 4; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 4; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 4; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 4; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 4; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 4; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 4; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 4; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 4; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 4; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 4; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 5; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 5; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 5; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 5; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 5; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 5; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 5; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 5; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 5; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 5; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 5; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 5; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 5; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 5; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 5; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 5; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 5; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 5; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 5; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 5; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 5; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 5; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 5; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 5; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 5; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 5; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 5; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 5; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 5; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 5; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 5; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 5; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 6; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 6; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 6; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 6; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 6; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 6; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 6; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 6; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 6; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 6; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 6; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 6; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 6; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 6; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 6; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 6; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 6; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 6; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 6; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 6; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 6; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 6; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 6; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 6; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 6; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 6; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 6; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 6; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 6; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 6; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 6; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 6; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 7; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 7; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 7; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 7; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 7; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 7; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 7; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 7; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 7; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 7; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 7; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 7; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 7; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 7; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 7; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 7; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 7; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 7; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 7; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 7; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 7; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 7; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 7; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 7; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 7; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 7; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 7; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 7; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 7; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 7; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 7; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 7; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 8; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 8; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 8; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 8; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 8; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 8; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 8; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 8; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 8; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 8; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 8; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 8; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 8; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 8; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 8; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 8; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 8; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 8; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 8; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 8; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 8; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 8; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 8; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 8; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 8; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 8; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 8; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 8; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 8; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 8; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 8; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 8; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 9; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 9; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 9; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 9; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 9; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 9; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 9; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 9; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 9; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 9; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 9; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 9; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 9; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 9; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 9; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 9; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 9; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 9; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 9; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 9; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 9; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 9; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 9; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 9; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 9; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 9; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 9; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 9; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 9; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 9; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 9; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 9; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 10; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 10; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 10; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 10; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 10; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 10; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 10; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 10; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 10; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 10; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 10; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 10; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 10; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 10; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 10; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 10; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 10; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 10; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 10; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 10; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 10; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 10; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 10; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 10; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 10; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 10; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 10; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 10; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 10; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 10; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 10; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 10; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 11; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 11; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 11; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 11; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 11; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 11; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 11; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 11; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 11; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 11; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 11; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 11; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 11; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 11; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 11; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 11; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 11; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 11; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 11; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 11; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 11; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 11; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 11; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 11; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 11; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 11; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 11; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 11; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 11; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 11; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 11; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 11; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 12; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 12; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 12; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 12; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 12; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 12; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 12; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 12; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 12; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 12; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 12; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 12; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 12; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 12; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 12; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 12; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 12; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 12; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 12; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 12; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 12; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 12; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 12; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 12; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 12; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 12; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 12; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 12; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 12; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 12; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 12; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 12; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 13; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 13; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 13; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 13; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 13; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 13; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 13; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 13; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 13; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 13; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 13; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 13; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 13; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 13; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 13; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 13; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 13; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 13; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 13; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 13; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 13; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 13; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 13; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 13; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 13; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 13; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 13; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 13; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 13; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 13; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 13; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 13; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 14; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 14; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 14; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 14; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 14; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 14; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 14; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 14; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 14; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 14; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 14; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 14; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 14; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 14; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 14; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 14; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 14; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 14; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 14; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 14; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 14; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 14; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 14; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 14; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 14; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 14; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 14; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 14; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 14; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 14; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 14; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 14; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 15; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 15; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 15; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 15; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 15; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 15; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 15; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 15; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 15; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 15; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 15; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 15; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 15; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 15; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 15; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 15; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 15; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 15; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 15; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 15; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 15; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 15; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 15; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 15; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 15; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 15; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 15; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 15; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 15; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 15; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 2; d1 <= 15; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 2; d1 <= 15; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 0; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 0; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 0; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 0; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 0; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 0; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 0; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 0; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 0; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 0; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 0; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 0; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 0; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 0; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 0; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 0; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 0; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 0; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 0; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 0; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 0; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 0; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 0; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 0; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 0; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 0; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 0; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 0; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 0; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 0; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 0; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 0; d0 <= 15; sel <= 1; // 
        #10 rst <= 0; sh_amt = 3; d1 <= 1; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 1; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 1; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 1; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 1; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 1; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 1; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 1; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 1; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 1; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 1; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 1; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 1; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 1; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 1; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 1; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 1; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 1; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 1; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 1; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 1; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 1; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 1; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 1; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 1; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 1; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 1; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 1; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 1; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 1; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 1; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 1; d0 <= 15; sel <= 1; // 
        #10 rst <= 0; sh_amt = 3; d1 <= 2; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 2; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 2; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 2; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 2; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 2; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 2; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 2; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 2; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 2; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 2; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 2; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 2; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 2; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 2; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 2; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 2; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 2; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 2; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 2; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 2; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 2; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 2; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 2; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 2; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 2; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 2; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 2; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 2; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 2; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 2; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 2; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 3; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 3; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 3; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 3; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 3; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 3; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 3; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 3; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 3; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 3; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 3; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 3; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 3; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 3; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 3; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 3; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 3; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 3; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 3; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 3; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 3; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 3; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 3; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 3; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 3; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 3; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 3; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 3; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 3; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 3; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 3; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 3; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 4; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 4; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 4; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 4; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 4; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 4; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 4; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 4; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 4; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 4; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 4; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 4; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 4; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 4; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 4; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 4; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 4; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 4; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 4; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 4; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 4; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 4; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 4; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 4; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 4; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 4; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 4; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 4; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 4; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 4; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 4; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 4; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 5; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 5; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 5; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 5; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 5; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 5; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 5; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 5; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 5; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 5; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 5; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 5; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 5; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 5; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 5; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 5; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 5; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 5; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 5; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 5; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 5; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 5; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 5; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 5; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 5; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 5; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 5; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 5; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 5; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 5; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 5; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 5; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 6; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 6; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 6; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 6; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 6; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 6; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 6; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 6; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 6; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 6; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 6; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 6; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 6; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 6; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 6; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 6; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 6; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 6; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 6; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 6; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 6; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 6; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 6; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 6; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 6; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 6; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 6; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 6; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 6; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 6; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 6; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 6; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 7; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 7; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 7; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 7; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 7; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 7; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 7; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 7; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 7; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 7; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 7; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 7; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 7; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 7; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 7; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 7; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 7; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 7; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 7; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 7; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 7; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 7; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 7; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 7; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 7; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 7; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 7; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 7; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 7; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 7; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 7; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 7; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 8; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 8; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 8; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 8; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 8; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 8; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 8; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 8; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 8; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 8; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 8; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 8; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 8; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 8; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 8; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 8; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 8; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 8; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 8; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 8; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 8; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 8; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 8; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 8; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 8; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 8; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 8; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 8; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 8; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 8; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 8; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 8; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 9; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 9; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 9; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 9; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 9; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 9; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 9; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 9; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 9; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 9; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 9; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 9; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 9; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 9; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 9; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 9; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 9; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 9; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 9; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 9; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 9; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 9; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 9; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 9; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 9; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 9; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 9; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 9; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 9; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 9; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 9; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 9; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 10; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 10; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 10; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 10; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 10; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 10; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 10; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 10; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 10; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 10; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 10; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 10; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 10; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 10; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 10; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 10; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 10; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 10; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 10; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 10; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 10; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 10; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 10; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 10; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 10; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 10; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 10; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 10; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 10; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 10; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 10; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 10; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 11; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 11; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 11; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 11; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 11; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 11; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 11; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 11; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 11; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 11; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 11; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 11; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 11; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 11; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 11; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 11; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 11; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 11; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 11; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 11; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 11; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 11; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 11; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 11; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 11; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 11; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 11; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 11; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 11; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 11; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 11; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 11; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 12; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 12; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 12; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 12; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 12; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 12; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 12; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 12; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 12; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 12; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 12; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 12; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 12; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 12; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 12; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 12; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 12; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 12; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 12; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 12; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 12; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 12; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 12; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 12; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 12; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 12; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 12; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 12; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 12; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 12; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 12; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 12; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 13; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 13; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 13; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 13; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 13; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 13; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 13; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 13; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 13; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 13; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 13; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 13; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 13; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 13; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 13; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 13; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 13; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 13; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 13; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 13; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 13; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 13; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 13; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 13; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 13; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 13; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 13; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 13; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 13; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 13; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 13; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 13; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 14; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 14; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 14; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 14; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 14; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 14; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 14; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 14; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 14; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 14; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 14; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 14; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 14; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 14; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 14; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 14; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 14; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 14; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 14; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 14; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 14; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 14; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 14; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 14; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 14; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 14; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 14; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 14; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 14; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 14; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 14; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 14; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 15; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 15; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 15; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 15; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 15; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 15; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 15; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 15; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 15; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 15; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 15; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 15; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 15; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 15; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 15; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 15; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 15; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 15; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 15; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 15; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 15; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 15; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 15; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 15; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 15; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 15; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 15; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 15; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 15; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 15; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 3; d1 <= 15; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 3; d1 <= 15; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 0; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 0; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 0; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 0; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 0; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 0; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 0; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 0; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 0; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 0; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 0; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 0; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 0; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 0; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 0; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 0; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 0; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 0; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 0; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 0; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 0; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 0; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 0; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 0; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 0; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 0; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 0; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 0; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 0; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 0; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 0; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 0; d0 <= 15; sel <= 1; // 
        #10 rst <= 0; sh_amt = 4; d1 <= 1; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 1; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 1; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 1; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 1; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 1; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 1; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 1; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 1; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 1; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 1; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 1; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 1; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 1; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 1; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 1; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 1; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 1; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 1; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 1; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 1; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 1; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 1; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 1; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 1; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 1; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 1; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 1; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 1; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 1; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 1; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 1; d0 <= 15; sel <= 1; // 
        #10 rst <= 0; sh_amt = 4; d1 <= 2; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 2; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 2; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 2; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 2; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 2; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 2; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 2; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 2; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 2; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 2; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 2; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 2; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 2; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 2; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 2; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 2; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 2; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 2; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 2; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 2; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 2; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 2; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 2; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 2; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 2; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 2; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 2; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 2; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 2; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 2; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 2; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 3; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 3; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 3; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 3; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 3; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 3; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 3; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 3; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 3; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 3; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 3; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 3; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 3; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 3; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 3; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 3; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 3; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 3; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 3; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 3; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 3; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 3; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 3; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 3; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 3; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 3; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 3; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 3; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 3; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 3; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 3; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 3; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 4; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 4; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 4; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 4; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 4; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 4; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 4; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 4; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 4; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 4; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 4; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 4; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 4; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 4; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 4; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 4; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 4; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 4; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 4; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 4; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 4; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 4; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 4; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 4; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 4; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 4; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 4; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 4; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 4; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 4; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 4; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 4; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 5; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 5; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 5; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 5; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 5; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 5; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 5; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 5; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 5; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 5; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 5; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 5; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 5; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 5; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 5; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 5; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 5; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 5; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 5; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 5; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 5; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 5; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 5; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 5; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 5; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 5; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 5; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 5; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 5; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 5; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 5; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 5; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 6; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 6; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 6; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 6; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 6; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 6; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 6; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 6; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 6; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 6; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 6; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 6; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 6; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 6; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 6; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 6; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 6; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 6; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 6; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 6; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 6; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 6; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 6; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 6; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 6; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 6; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 6; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 6; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 6; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 6; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 6; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 6; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 7; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 7; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 7; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 7; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 7; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 7; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 7; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 7; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 7; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 7; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 7; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 7; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 7; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 7; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 7; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 7; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 7; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 7; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 7; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 7; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 7; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 7; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 7; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 7; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 7; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 7; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 7; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 7; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 7; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 7; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 7; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 7; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 8; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 8; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 8; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 8; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 8; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 8; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 8; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 8; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 8; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 8; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 8; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 8; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 8; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 8; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 8; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 8; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 8; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 8; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 8; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 8; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 8; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 8; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 8; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 8; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 8; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 8; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 8; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 8; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 8; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 8; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 8; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 8; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 9; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 9; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 9; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 9; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 9; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 9; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 9; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 9; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 9; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 9; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 9; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 9; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 9; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 9; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 9; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 9; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 9; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 9; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 9; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 9; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 9; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 9; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 9; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 9; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 9; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 9; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 9; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 9; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 9; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 9; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 9; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 9; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 10; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 10; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 10; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 10; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 10; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 10; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 10; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 10; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 10; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 10; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 10; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 10; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 10; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 10; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 10; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 10; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 10; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 10; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 10; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 10; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 10; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 10; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 10; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 10; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 10; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 10; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 10; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 10; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 10; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 10; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 10; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 10; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 11; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 11; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 11; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 11; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 11; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 11; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 11; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 11; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 11; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 11; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 11; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 11; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 11; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 11; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 11; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 11; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 11; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 11; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 11; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 11; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 11; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 11; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 11; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 11; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 11; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 11; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 11; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 11; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 11; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 11; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 11; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 11; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 12; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 12; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 12; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 12; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 12; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 12; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 12; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 12; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 12; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 12; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 12; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 12; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 12; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 12; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 12; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 12; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 12; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 12; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 12; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 12; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 12; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 12; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 12; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 12; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 12; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 12; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 12; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 12; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 12; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 12; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 12; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 12; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 13; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 13; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 13; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 13; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 13; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 13; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 13; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 13; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 13; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 13; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 13; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 13; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 13; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 13; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 13; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 13; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 13; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 13; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 13; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 13; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 13; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 13; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 13; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 13; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 13; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 13; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 13; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 13; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 13; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 13; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 13; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 13; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 14; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 14; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 14; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 14; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 14; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 14; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 14; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 14; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 14; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 14; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 14; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 14; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 14; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 14; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 14; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 14; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 14; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 14; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 14; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 14; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 14; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 14; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 14; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 14; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 14; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 14; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 14; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 14; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 14; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 14; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 14; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 14; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 15; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 15; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 15; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 15; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 15; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 15; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 15; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 15; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 15; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 15; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 15; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 15; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 15; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 15; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 15; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 15; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 15; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 15; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 15; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 15; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 15; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 15; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 15; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 15; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 15; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 15; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 15; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 15; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 15; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 15; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 4; d1 <= 15; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 4; d1 <= 15; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 0; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 0; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 0; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 0; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 0; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 0; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 0; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 0; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 0; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 0; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 0; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 0; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 0; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 0; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 0; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 0; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 0; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 0; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 0; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 0; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 0; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 0; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 0; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 0; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 0; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 0; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 0; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 0; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 0; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 0; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 0; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 0; d0 <= 15; sel <= 1; // 
        #10 rst <= 0; sh_amt = 5; d1 <= 1; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 1; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 1; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 1; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 1; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 1; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 1; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 1; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 1; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 1; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 1; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 1; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 1; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 1; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 1; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 1; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 1; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 1; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 1; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 1; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 1; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 1; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 1; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 1; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 1; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 1; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 1; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 1; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 1; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 1; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 1; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 1; d0 <= 15; sel <= 1; // 
        #10 rst <= 0; sh_amt = 5; d1 <= 2; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 2; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 2; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 2; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 2; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 2; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 2; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 2; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 2; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 2; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 2; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 2; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 2; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 2; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 2; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 2; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 2; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 2; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 2; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 2; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 2; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 2; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 2; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 2; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 2; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 2; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 2; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 2; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 2; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 2; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 2; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 2; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 3; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 3; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 3; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 3; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 3; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 3; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 3; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 3; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 3; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 3; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 3; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 3; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 3; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 3; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 3; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 3; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 3; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 3; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 3; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 3; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 3; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 3; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 3; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 3; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 3; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 3; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 3; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 3; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 3; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 3; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 3; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 3; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 4; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 4; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 4; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 4; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 4; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 4; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 4; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 4; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 4; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 4; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 4; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 4; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 4; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 4; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 4; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 4; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 4; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 4; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 4; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 4; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 4; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 4; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 4; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 4; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 4; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 4; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 4; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 4; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 4; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 4; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 4; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 4; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 5; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 5; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 5; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 5; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 5; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 5; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 5; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 5; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 5; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 5; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 5; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 5; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 5; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 5; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 5; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 5; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 5; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 5; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 5; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 5; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 5; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 5; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 5; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 5; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 5; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 5; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 5; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 5; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 5; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 5; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 5; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 5; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 6; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 6; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 6; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 6; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 6; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 6; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 6; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 6; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 6; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 6; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 6; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 6; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 6; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 6; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 6; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 6; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 6; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 6; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 6; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 6; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 6; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 6; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 6; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 6; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 6; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 6; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 6; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 6; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 6; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 6; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 6; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 6; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 7; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 7; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 7; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 7; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 7; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 7; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 7; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 7; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 7; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 7; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 7; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 7; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 7; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 7; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 7; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 7; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 7; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 7; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 7; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 7; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 7; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 7; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 7; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 7; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 7; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 7; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 7; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 7; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 7; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 7; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 7; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 7; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 8; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 8; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 8; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 8; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 8; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 8; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 8; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 8; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 8; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 8; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 8; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 8; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 8; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 8; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 8; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 8; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 8; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 8; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 8; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 8; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 8; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 8; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 8; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 8; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 8; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 8; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 8; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 8; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 8; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 8; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 8; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 8; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 9; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 9; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 9; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 9; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 9; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 9; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 9; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 9; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 9; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 9; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 9; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 9; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 9; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 9; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 9; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 9; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 9; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 9; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 9; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 9; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 9; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 9; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 9; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 9; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 9; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 9; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 9; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 9; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 9; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 9; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 9; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 9; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 10; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 10; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 10; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 10; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 10; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 10; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 10; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 10; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 10; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 10; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 10; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 10; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 10; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 10; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 10; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 10; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 10; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 10; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 10; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 10; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 10; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 10; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 10; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 10; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 10; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 10; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 10; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 10; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 10; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 10; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 10; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 10; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 11; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 11; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 11; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 11; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 11; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 11; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 11; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 11; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 11; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 11; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 11; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 11; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 11; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 11; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 11; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 11; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 11; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 11; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 11; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 11; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 11; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 11; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 11; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 11; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 11; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 11; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 11; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 11; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 11; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 11; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 11; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 11; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 12; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 12; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 12; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 12; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 12; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 12; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 12; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 12; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 12; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 12; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 12; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 12; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 12; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 12; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 12; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 12; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 12; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 12; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 12; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 12; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 12; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 12; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 12; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 12; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 12; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 12; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 12; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 12; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 12; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 12; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 12; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 12; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 13; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 13; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 13; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 13; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 13; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 13; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 13; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 13; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 13; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 13; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 13; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 13; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 13; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 13; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 13; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 13; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 13; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 13; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 13; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 13; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 13; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 13; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 13; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 13; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 13; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 13; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 13; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 13; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 13; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 13; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 13; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 13; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 14; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 14; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 14; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 14; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 14; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 14; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 14; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 14; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 14; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 14; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 14; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 14; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 14; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 14; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 14; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 14; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 14; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 14; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 14; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 14; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 14; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 14; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 14; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 14; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 14; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 14; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 14; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 14; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 14; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 14; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 14; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 14; d0 <= 15; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 15; d0 <= 0; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 15; d0 <= 0; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 15; d0 <= 1; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 15; d0 <= 1; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 15; d0 <= 2; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 15; d0 <= 2; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 15; d0 <= 3; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 15; d0 <= 3; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 15; d0 <= 4; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 15; d0 <= 4; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 15; d0 <= 5; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 15; d0 <= 5; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 15; d0 <= 6; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 15; d0 <= 6; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 15; d0 <= 7; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 15; d0 <= 7; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 15; d0 <= 8; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 15; d0 <= 8; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 15; d0 <= 9; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 15; d0 <= 9; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 15; d0 <= 10; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 15; d0 <= 10; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 15; d0 <= 11; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 15; d0 <= 11; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 15; d0 <= 12; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 15; d0 <= 12; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 15; d0 <= 13; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 15; d0 <= 13; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 15; d0 <= 14; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 15; d0 <= 14; sel <= 1; 
        #10 rst <= 0; sh_amt = 5; d1 <= 15; d0 <= 15; sel <= 0; 
        #10 rst <= 0; sh_amt = 5; d1 <= 15; d0 <= 15; sel <= 1; 
    end
    
    always begin
        #5 clk <= ~clk;
    end
endmodule
